`timescale 1 ns / 1 ps



module mnist_nn_tb();


reg clk,reset;
reg inp_ready;
reg [15:0] inp_data;

wire [15:0] w_0, w_1;

wire [9:0] inp_count;



wire [7:0] n0_out, n1_out;

wire n1_ready,n0_ready;



initial begin
	clk = 1'b1;
	forever #1 clk = ~clk;
end


initial
#2000 $stop;

//initial
//begin
//reset = 1'b1;
//#1 reset = 1'b0;
//end


mnist_nn mnist_dut(.clk(clk),
				   .reset(reset),
				   .inp_rdy(inp_ready),
				   .inp_data(inp_data),
				   
				   .inp_count(inp_count),
				   .weight_value_0(w_0),
				   .weight_value_1(w_1),
				   .n0_out(n0_out),
				   .n1_out(n1_out),
				   .n0_ready(n0_ready),
				   .n1_ready(n1_ready)
				   
				   );


initial begin
        
        reset = 1;
        inp_ready = 0;
        inp_data = 0;


        #5 reset = 0; 

        #5;
		
		inp_ready = 1;
		
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h000b; #2
		inp_data = 16'h0097; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00cb; #2
		inp_data = 16'h001f; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0025; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h006b; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0015; #2
		inp_data = 16'h00c6; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h006b; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h006e; #2
		inp_data = 16'h00bf; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00aa; #2
		inp_data = 16'h006d; #2
		inp_data = 16'h003e; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00dd; #2
		inp_data = 16'h0033; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00b7; #2
		inp_data = 16'h0100; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00eb; #2
		inp_data = 16'h00df; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h003f; #2
		inp_data = 16'h00de; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0094; #2
		inp_data = 16'h004d; #2
		inp_data = 16'h003e; #2
		inp_data = 16'h0081; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0069; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0020; #2
		inp_data = 16'h00e8; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00dd; #2
		inp_data = 16'h008a; #2
		inp_data = 16'h000a; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h001f; #2
		inp_data = 16'h00e7; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00f4; #2
		inp_data = 16'h0071; #2
		inp_data = 16'h0005; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0025; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00bd; #2
		inp_data = 16'h0014; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h006d; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0023; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0025; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00ca; #2
		inp_data = 16'h001e; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h001f; #2
		inp_data = 16'h00c9; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0023; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0025; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0020; #2
		inp_data = 16'h00cb; #2
		inp_data = 16'h0100; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00a5; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h008d; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h006d; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0023; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00da; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0015; #2
		inp_data = 16'h003f; #2
		inp_data = 16'h00e8; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00e7; #2
		inp_data = 16'h001e; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00da; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0091; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00de; #2
		inp_data = 16'h003d; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00da; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00b7; #2
		inp_data = 16'h00de; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00b5; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h00db; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h0049; #2
		inp_data = 16'h0049; #2
		inp_data = 16'h00e5; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h0100; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0071; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h0094; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h001f; #2
		inp_data = 16'h00e7; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00e7; #2
		inp_data = 16'h00be; #2
		inp_data = 16'h0023; #2
		inp_data = 16'h000a; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h003e; #2
		inp_data = 16'h008f; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00fe; #2
		inp_data = 16'h006b; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0048; #2
		inp_data = 16'h00af; #2
		inp_data = 16'h00fc; #2
		inp_data = 16'h00ae; #2
		inp_data = 16'h0047; #2
		inp_data = 16'h0048; #2
		inp_data = 16'h001e; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		inp_data = 16'h0000; #2
		
		inp_ready = 0;


end





				   
				   
endmodule