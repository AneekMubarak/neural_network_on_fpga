`timescale 1 ns / 1 ps


module neuron_tb();



	reg clk,reset,inp_ready;

	reg signed [15:0] inp_data, weight, bias;

	wire out_ready;


	wire [31:0] product_q16_16, acc_final, acc ;
	 
	wire [9:0] count;
	
	wire [11:0] sig_addr;
	
	wire [7:0] sig_out;
	
	wire sig_ready;
	
	
	



	neuron neuron_dut(
					.clk(clk),
					.reset(reset),
					.inp_data(inp_data),
					.weight(weight),
					.bias(bias),
					.out_ready(out_ready),
					.acc_final(acc_final),
					.product_q16_16(product_q16_16),
					.acc(acc),
					.count(count),
					.inp_ready(inp_ready),
					.sigmoid_out(sig_out),
					.sigmoid_address(sig_addr),
					.sigmoid_ready(sig_ready)
					);
 
	initial
	#2000 $stop; 
	 
	initial 
		begin
			clk = 1'b1;
			forever #1 clk = ~clk;
		end
	
	
 
// test 1: check product calculation
// test 2: check output and format for mathematical accuracy
// test 3: check out_ready_signal
    initial begin
        
        reset = 1;
        inp_ready = 0;
        inp_data = 0;
        weight = 0;
        bias = 0;

        #5 reset = 0; 

        #5;
		
		bias = 16'hff4b;
		inp_ready = 1;


        // inp_data = 1.5 (in Q8.8) = 16'h0180
        // weight = -2.0 (Q8.8) = 16'hfe00
        // inp_data = 16'h080; // 1.5
        // weight = 16'hFE00;   // -2.0
		

		// #2 //full clk cyclr
		// inp_data = 16'h00ff;
		// weight   = 16'hffff;
		
		
		// #2 
		// inp_data = 16'h0012;
		// weight   = 16'hffff;
		
		
		// #2 
		// inp_data = 16'h0000;
		// weight   = 16'h0000;
		        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'hfff4; #2;
        inp_data = 16'h0000; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hffde; #2;
        inp_data = 16'h0000; weight = 16'hffd5; #2;
        inp_data = 16'h0000; weight = 16'hffe5; #2;
        inp_data = 16'h0000; weight = 16'hffdd; #2;
        inp_data = 16'h0000; weight = 16'hffe6; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'hfff4; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0010; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h000b; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hffde; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hffe3; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0032; weight = 16'h0024; #2;
        inp_data = 16'h00e1; weight = 16'h0014; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0025; #2;
        inp_data = 16'h0000; weight = 16'h003f; #2;
        inp_data = 16'h0000; weight = 16'h0025; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'h003e; #2;
        inp_data = 16'h0000; weight = 16'h003f; #2;
        inp_data = 16'h0046; weight = 16'h0011; #2;
        inp_data = 16'h001d; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hffd8; #2;
        inp_data = 16'h0000; weight = 16'hffdf; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'hffe3; #2;
        inp_data = 16'h0079; weight = 16'h000e; #2;
        inp_data = 16'h00e8; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'h002b; #2;
        inp_data = 16'h0000; weight = 16'h0023; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h001f; #2;
        inp_data = 16'h0000; weight = 16'h002f; #2;
        inp_data = 16'h0000; weight = 16'h0042; #2;
        inp_data = 16'h0095; weight = 16'h0021; #2;
        inp_data = 16'h00a9; weight = 16'h0018; #2;
        inp_data = 16'h0000; weight = 16'h003d; #2;
        inp_data = 16'h0000; weight = 16'h0038; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hffcb; #2;
        inp_data = 16'h0000; weight = 16'hffd8; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hffd6; #2;
        inp_data = 16'h0004; weight = 16'hfffe; #2;
        inp_data = 16'h00c4; weight = 16'h000d; #2;
        inp_data = 16'h00e8; weight = 16'h000e; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h001f; #2;
        inp_data = 16'h0000; weight = 16'h0019; #2;
        inp_data = 16'h0000; weight = 16'h000e; #2;
        inp_data = 16'h0000; weight = 16'h000e; #2;
        inp_data = 16'h0000; weight = 16'h003f; #2;
        inp_data = 16'h0000; weight = 16'h003c; #2;
        inp_data = 16'h0060; weight = 16'h002c; #2;
        inp_data = 16'h00d3; weight = 16'h0009; #2;
        inp_data = 16'h000b; weight = 16'h000f; #2;
        inp_data = 16'h0000; weight = 16'h0026; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'hffe2; #2;
        inp_data = 16'h0000; weight = 16'hffd1; #2;
        inp_data = 16'h0000; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hffe9; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0045; weight = 16'h001b; #2;
        inp_data = 16'h00fd; weight = 16'h0011; #2;
        inp_data = 16'h0087; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0017; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h002a; #2;
        inp_data = 16'h0000; weight = 16'h003b; #2;
        inp_data = 16'h0000; weight = 16'h006d; #2;
        inp_data = 16'h0000; weight = 16'h0048; #2;
        inp_data = 16'h0000; weight = 16'h0035; #2;
        inp_data = 16'h0072; weight = 16'h000f; #2;
        inp_data = 16'h00fd; weight = 16'h0017; #2;
        inp_data = 16'h0015; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'h002a; #2;
        inp_data = 16'h0000; weight = 16'h0059; #2;
        inp_data = 16'h0000; weight = 16'h000b; #2;
        inp_data = 16'h0000; weight = 16'hffd0; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hffee; #2;
        inp_data = 16'h0000; weight = 16'hffe5; #2;
        inp_data = 16'h002d; weight = 16'hffe6; #2;
        inp_data = 16'h00ed; weight = 16'hfffd; #2;
        inp_data = 16'h00da; weight = 16'h001c; #2;
        inp_data = 16'h000c; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h003c; #2;
        inp_data = 16'h0000; weight = 16'h0012; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'h002e; #2;
        inp_data = 16'h0000; weight = 16'h0045; #2;
        inp_data = 16'h0000; weight = 16'h004a; #2;
        inp_data = 16'h00c1; weight = 16'h0036; #2;
        inp_data = 16'h00fd; weight = 16'h0022; #2;
        inp_data = 16'h0015; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h001a; #2;
        inp_data = 16'h0000; weight = 16'h0060; #2;
        inp_data = 16'h0000; weight = 16'h0028; #2;
        inp_data = 16'h0000; weight = 16'hffcd; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hffe3; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h00a9; weight = 16'hfff2; #2;
        inp_data = 16'h00f8; weight = 16'h0007; #2;
        inp_data = 16'h0035; weight = 16'hffe4; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0013; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hffd9; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h004c; #2;
        inp_data = 16'h0012; weight = 16'h0043; #2;
        inp_data = 16'h0100; weight = 16'h0017; #2;
        inp_data = 16'h00fe; weight = 16'h0025; #2;
        inp_data = 16'h0015; weight = 16'h0012; #2;
        inp_data = 16'h0000; weight = 16'h0031; #2;
        inp_data = 16'h0000; weight = 16'h0067; #2;
        inp_data = 16'h0000; weight = 16'h0038; #2;
        inp_data = 16'h0000; weight = 16'hffd3; #2;
        inp_data = 16'h0000; weight = 16'hffe6; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hffde; #2;
        inp_data = 16'h0000; weight = 16'hffe9; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0054; weight = 16'h0005; #2;
        inp_data = 16'h00f3; weight = 16'h0002; #2;
        inp_data = 16'h00d4; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hffdd; #2;
        inp_data = 16'h0000; weight = 16'hfff4; #2;
        inp_data = 16'h0000; weight = 16'hffab; #2;
        inp_data = 16'h0000; weight = 16'hff71; #2;
        inp_data = 16'h0000; weight = 16'hff7b; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h008e; weight = 16'hfff0; #2;
        inp_data = 16'h00fe; weight = 16'h000c; #2;
        inp_data = 16'h00be; weight = 16'h002b; #2;
        inp_data = 16'h0005; weight = 16'h003c; #2;
        inp_data = 16'h0000; weight = 16'h0042; #2;
        inp_data = 16'h0000; weight = 16'h0055; #2;
        inp_data = 16'h0000; weight = 16'h0043; #2;
        inp_data = 16'h0000; weight = 16'hffd9; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hffe9; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0023; #2;
        inp_data = 16'h00aa; weight = 16'h0009; #2;
        inp_data = 16'h00fd; weight = 16'hfff3; #2;
        inp_data = 16'h006a; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'h000b; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0011; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'hff79; #2;
        inp_data = 16'h0000; weight = 16'hff43; #2;
        inp_data = 16'h0000; weight = 16'hff64; #2;
        inp_data = 16'h0020; weight = 16'hffda; #2;
        inp_data = 16'h00e9; weight = 16'hfff2; #2;
        inp_data = 16'h00fb; weight = 16'h000f; #2;
        inp_data = 16'h0042; weight = 16'h0013; #2;
        inp_data = 16'h0000; weight = 16'h001f; #2;
        inp_data = 16'h0000; weight = 16'h0044; #2;
        inp_data = 16'h0000; weight = 16'h006a; #2;
        inp_data = 16'h0000; weight = 16'h0063; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h000f; weight = 16'h0045; #2;
        inp_data = 16'h00e2; weight = 16'h0040; #2;
        inp_data = 16'h00fd; weight = 16'h0019; #2;
        inp_data = 16'h0000; weight = 16'h0016; #2;
        inp_data = 16'h0000; weight = 16'h0024; #2;
        inp_data = 16'h0000; weight = 16'h0013; #2;
        inp_data = 16'h0000; weight = 16'h0014; #2;
        inp_data = 16'h0000; weight = 16'hffa7; #2;
        inp_data = 16'h0000; weight = 16'hff63; #2;
        inp_data = 16'h0000; weight = 16'hff31; #2;
        inp_data = 16'h0000; weight = 16'hff6d; #2;
        inp_data = 16'h0087; weight = 16'hffc4; #2;
        inp_data = 16'h00fd; weight = 16'hfffa; #2;
        inp_data = 16'h00d4; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'hffcb; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0036; #2;
        inp_data = 16'h0000; weight = 16'h0062; #2;
        inp_data = 16'h0000; weight = 16'h005f; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'h0039; #2;
        inp_data = 16'h0016; weight = 16'h003a; #2;
        inp_data = 16'h00fd; weight = 16'h0056; #2;
        inp_data = 16'h00a5; weight = 16'h0035; #2;
        inp_data = 16'h0000; weight = 16'h003a; #2;
        inp_data = 16'h0000; weight = 16'h0023; #2;
        inp_data = 16'h0000; weight = 16'h0031; #2;
        inp_data = 16'h0000; weight = 16'h0020; #2;
        inp_data = 16'h0000; weight = 16'hffb6; #2;
        inp_data = 16'h0000; weight = 16'hff4d; #2;
        inp_data = 16'h0000; weight = 16'hff4d; #2;
        inp_data = 16'h0000; weight = 16'hff57; #2;
        inp_data = 16'h00aa; weight = 16'hffd8; #2;
        inp_data = 16'h00fd; weight = 16'hffed; #2;
        inp_data = 16'h00a8; weight = 16'hffdc; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0022; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'h0058; #2;
        inp_data = 16'h0000; weight = 16'h0054; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0013; #2;
        inp_data = 16'h0000; weight = 16'h0050; #2;
        inp_data = 16'h0009; weight = 16'h0015; #2;
        inp_data = 16'h00cd; weight = 16'h004d; #2;
        inp_data = 16'h00d2; weight = 16'h003e; #2;
        inp_data = 16'h0012; weight = 16'h003d; #2;
        inp_data = 16'h0000; weight = 16'h0045; #2;
        inp_data = 16'h0000; weight = 16'h0014; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'hff7f; #2;
        inp_data = 16'h0000; weight = 16'hff2a; #2;
        inp_data = 16'h0000; weight = 16'hff61; #2;
        inp_data = 16'h0016; weight = 16'hff87; #2;
        inp_data = 16'h00fe; weight = 16'hffcb; #2;
        inp_data = 16'h00fe; weight = 16'hfff5; #2;
        inp_data = 16'h006b; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'h0023; #2;
        inp_data = 16'h0000; weight = 16'h0019; #2;
        inp_data = 16'h0000; weight = 16'h002a; #2;
        inp_data = 16'h0000; weight = 16'h0058; #2;
        inp_data = 16'h0000; weight = 16'h0048; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hffec; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'h0056; #2;
        inp_data = 16'h0000; weight = 16'h0039; #2;
        inp_data = 16'h00aa; weight = 16'h003e; #2;
        inp_data = 16'h00fd; weight = 16'h0048; #2;
        inp_data = 16'h00c8; weight = 16'h0048; #2;
        inp_data = 16'h0055; weight = 16'h003e; #2;
        inp_data = 16'h0055; weight = 16'h0017; #2;
        inp_data = 16'h0055; weight = 16'hffb9; #2;
        inp_data = 16'h0055; weight = 16'hff41; #2;
        inp_data = 16'h0082; weight = 16'hff4e; #2;
        inp_data = 16'h00a5; weight = 16'hff8d; #2;
        inp_data = 16'h00c4; weight = 16'hffc4; #2;
        inp_data = 16'h00fd; weight = 16'hfff8; #2;
        inp_data = 16'h00fd; weight = 16'h0004; #2;
        inp_data = 16'h006a; weight = 16'h000b; #2;
        inp_data = 16'h0000; weight = 16'h0034; #2;
        inp_data = 16'h0000; weight = 16'h0021; #2;
        inp_data = 16'h0000; weight = 16'h002d; #2;
        inp_data = 16'h0000; weight = 16'h0037; #2;
        inp_data = 16'h0000; weight = 16'h0018; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0012; #2;
        inp_data = 16'h0000; weight = 16'h0042; #2;
        inp_data = 16'h0000; weight = 16'h0039; #2;
        inp_data = 16'h0029; weight = 16'h002f; #2;
        inp_data = 16'h00ab; weight = 16'h001c; #2;
        inp_data = 16'h00f6; weight = 16'h0043; #2;
        inp_data = 16'h00fd; weight = 16'h0067; #2;
        inp_data = 16'h00fd; weight = 16'h0020; #2;
        inp_data = 16'h00fd; weight = 16'hffd0; #2;
        inp_data = 16'h00fd; weight = 16'hff63; #2;
        inp_data = 16'h00e9; weight = 16'hff68; #2;
        inp_data = 16'h00e8; weight = 16'hffb0; #2;
        inp_data = 16'h00fc; weight = 16'hfff2; #2;
        inp_data = 16'h00fd; weight = 16'h001b; #2;
        inp_data = 16'h00fd; weight = 16'h0004; #2;
        inp_data = 16'h0009; weight = 16'h0012; #2;
        inp_data = 16'h0000; weight = 16'h001e; #2;
        inp_data = 16'h0000; weight = 16'h000e; #2;
        inp_data = 16'h0000; weight = 16'h0029; #2;
        inp_data = 16'h0000; weight = 16'h0014; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0021; #2;
        inp_data = 16'h0000; weight = 16'h0028; #2;
        inp_data = 16'h0000; weight = 16'h0020; #2;
        inp_data = 16'h0000; weight = 16'h003b; #2;
        inp_data = 16'h0031; weight = 16'h003f; #2;
        inp_data = 16'h0054; weight = 16'h0058; #2;
        inp_data = 16'h0054; weight = 16'h0017; #2;
        inp_data = 16'h0054; weight = 16'hffc2; #2;
        inp_data = 16'h0054; weight = 16'hff69; #2;
        inp_data = 16'h0000; weight = 16'hff92; #2;
        inp_data = 16'h0000; weight = 16'hffd3; #2;
        inp_data = 16'h00a2; weight = 16'hfff2; #2;
        inp_data = 16'h00fd; weight = 16'h0005; #2;
        inp_data = 16'h00fd; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0032; #2;
        inp_data = 16'h0000; weight = 16'h0012; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hffee; #2;
        inp_data = 16'h0000; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'h0021; #2;
        inp_data = 16'h0000; weight = 16'h0030; #2;
        inp_data = 16'h0000; weight = 16'h003f; #2;
        inp_data = 16'h0000; weight = 16'h0034; #2;
        inp_data = 16'h0000; weight = 16'h0029; #2;
        inp_data = 16'h0000; weight = 16'h004f; #2;
        inp_data = 16'h0000; weight = 16'h0052; #2;
        inp_data = 16'h0000; weight = 16'h0031; #2;
        inp_data = 16'h0000; weight = 16'hffd6; #2;
        inp_data = 16'h0000; weight = 16'hffcd; #2;
        inp_data = 16'h0000; weight = 16'hffdf; #2;
        inp_data = 16'h007f; weight = 16'hffec; #2;
        inp_data = 16'h00fd; weight = 16'h0006; #2;
        inp_data = 16'h00fd; weight = 16'h0000; #2;
        inp_data = 16'h002d; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0018; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h000b; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'h002e; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'h001c; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'h0027; #2;
        inp_data = 16'h0000; weight = 16'h005c; #2;
        inp_data = 16'h0000; weight = 16'h006c; #2;
        inp_data = 16'h0000; weight = 16'h0065; #2;
        inp_data = 16'h0000; weight = 16'h0030; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0081; weight = 16'hffef; #2;
        inp_data = 16'h00fe; weight = 16'h0003; #2;
        inp_data = 16'h00fe; weight = 16'hffe0; #2;
        inp_data = 16'h0000; weight = 16'hffd6; #2;
        inp_data = 16'h0000; weight = 16'hffea; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0014; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfff1; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'h001c; #2;
        inp_data = 16'h0000; weight = 16'h0022; #2;
        inp_data = 16'h0000; weight = 16'h001c; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h000c; #2;
        inp_data = 16'h0000; weight = 16'h003d; #2;
        inp_data = 16'h0000; weight = 16'h0057; #2;
        inp_data = 16'h0000; weight = 16'h0047; #2;
        inp_data = 16'h0000; weight = 16'h001d; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h007f; weight = 16'hfffc; #2;
        inp_data = 16'h00fd; weight = 16'hffc9; #2;
        inp_data = 16'h00fd; weight = 16'hffcb; #2;
        inp_data = 16'h0000; weight = 16'hffc6; #2;
        inp_data = 16'h0000; weight = 16'hffee; #2;
        inp_data = 16'h0000; weight = 16'h000a; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hffec; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hffd2; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0010; #2;
        inp_data = 16'h0000; weight = 16'h000e; #2;
        inp_data = 16'h0000; weight = 16'h0028; #2;
        inp_data = 16'h0000; weight = 16'h001f; #2;
        inp_data = 16'h0000; weight = 16'h0024; #2;
        inp_data = 16'h0000; weight = 16'h0031; #2;
        inp_data = 16'h0000; weight = 16'h0029; #2;
        inp_data = 16'h0000; weight = 16'h0066; #2;
        inp_data = 16'h0000; weight = 16'h002d; #2;
        inp_data = 16'h0000; weight = 16'h001c; #2;
        inp_data = 16'h0088; weight = 16'h0007; #2;
        inp_data = 16'h00fd; weight = 16'h0006; #2;
        inp_data = 16'h00f5; weight = 16'hffe1; #2;
        inp_data = 16'h0000; weight = 16'hffe2; #2;
        inp_data = 16'h0000; weight = 16'hffd6; #2;
        inp_data = 16'h0000; weight = 16'hffe5; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hffdd; #2;
        inp_data = 16'h0000; weight = 16'hffdc; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'h001d; #2;
        inp_data = 16'h0000; weight = 16'h0037; #2;
        inp_data = 16'h0000; weight = 16'h0056; #2;
        inp_data = 16'h0000; weight = 16'h005e; #2;
        inp_data = 16'h0000; weight = 16'h0045; #2;
        inp_data = 16'h0000; weight = 16'h0045; #2;
        inp_data = 16'h0000; weight = 16'h0039; #2;
        inp_data = 16'h0000; weight = 16'h0028; #2;
        inp_data = 16'h00e9; weight = 16'hfffb; #2;
        inp_data = 16'h00ed; weight = 16'h0006; #2;
        inp_data = 16'h006f; weight = 16'hffc4; #2;
        inp_data = 16'h0000; weight = 16'hffbe; #2;
        inp_data = 16'h0000; weight = 16'hffc0; #2;
        inp_data = 16'h0000; weight = 16'hffdd; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0007; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'hffe1; #2;
        inp_data = 16'h0000; weight = 16'hffdc; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hffee; #2;
        inp_data = 16'h0000; weight = 16'hfff4; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0025; #2;
        inp_data = 16'h0000; weight = 16'h0030; #2;
        inp_data = 16'h0000; weight = 16'h0013; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h00b4; weight = 16'hffde; #2;
        inp_data = 16'h0042; weight = 16'hffd9; #2;
        inp_data = 16'h0000; weight = 16'hffc9; #2;
        inp_data = 16'h0000; weight = 16'hffca; #2;
        inp_data = 16'h0000; weight = 16'hffca; #2;
        inp_data = 16'h0000; weight = 16'hffe4; #2;
        inp_data = 16'h0000; weight = 16'hfff2; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfff5; #2;
        inp_data = 16'h0000; weight = 16'hfff6; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hffd1; #2;
        inp_data = 16'h0000; weight = 16'hffc8; #2;
        inp_data = 16'h0000; weight = 16'hffaf; #2;
        inp_data = 16'h0000; weight = 16'hffb6; #2;
        inp_data = 16'h0000; weight = 16'hffad; #2;
        inp_data = 16'h0000; weight = 16'hffad; #2;
        inp_data = 16'h0000; weight = 16'hffb9; #2;
        inp_data = 16'h0000; weight = 16'hffbf; #2;
        inp_data = 16'h0000; weight = 16'hffce; #2;
        inp_data = 16'h0000; weight = 16'hffc2; #2;
        inp_data = 16'h0000; weight = 16'hffcf; #2;
        inp_data = 16'h0000; weight = 16'hffdf; #2;
        inp_data = 16'h0000; weight = 16'hffdf; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0006; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff8; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfff0; #2;
        inp_data = 16'h0000; weight = 16'hffe7; #2;
        inp_data = 16'h0000; weight = 16'hfff3; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hffef; #2;
        inp_data = 16'h0000; weight = 16'hffeb; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hffed; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff4; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'h0000; #2;
        inp_data = 16'h0000; weight = 16'h0004; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'h0009; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfffa; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'h0005; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'hfff7; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'h0008; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hfffb; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'hfff9; #2;
        inp_data = 16'h0000; weight = 16'hffff; #2;
        inp_data = 16'h0000; weight = 16'hfffd; #2;
        inp_data = 16'h0000; weight = 16'hfffe; #2;
        inp_data = 16'h0000; weight = 16'h0001; #2;
        inp_data = 16'h0000; weight = 16'hfffc; #2;
        inp_data = 16'h0000; weight = 16'h0002; #2;
        inp_data = 16'h0000; weight = 16'h0003; #2;


 
    end

endmodule








// test 2: check output and format for mathematical accuracy

// test 3: check out_ready_signal